module Datapath #(
    parameter N = 64
)(
    input  logic       clk, rst,
    input  logic       regWriteEnable,
    input  logic       memWriteEnable,
    input  logic       ALU_srcB_sel, result_src_sel, pc_src_sel
);



endmodule
